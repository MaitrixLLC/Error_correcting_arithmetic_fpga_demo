// q_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module q_sys (
		input  wire        clk_clk,                                      //                                   clk.clk
		input  wire [9:0]  in_fifo_used_external_connection_export,      //      in_fifo_used_external_connection.export
		input  wire [31:0] in_port_data_external_connection_export,      //      in_port_data_external_connection.export
		input  wire [19:0] in_port_dig_error_external_connection_export, // in_port_dig_error_external_connection.export
		input  wire [2:0]  in_port_ec_flags_external_connection_export,  //  in_port_ec_flags_external_connection.export
		input  wire [15:0] in_port_freq_cnt_external_connection_export,  //  in_port_freq_cnt_external_connection.export
		output wire [9:0]  out_port_batnum_external_connection_export,   //   out_port_batnum_external_connection.export
		output wire [7:0]  out_port_ctrl_external_connection_export,     //     out_port_ctrl_external_connection.export
		output wire [10:0] out_port_lut_adr_external_connection_export,  //  out_port_lut_adr_external_connection.export
		output wire [31:0] out_port_lut_data_external_connection_export, // out_port_lut_data_external_connection.export
		output wire [9:0]  out_port_prodnum_external_connection_export,  //  out_port_prodnum_external_connection.export
		input  wire        reset_reset_n,                                //                                 reset.reset_n
		input  wire        uart_0_external_connection_rxd,               //            uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd                //                                      .txd
	);

	wire         pll_0_50_outclk0_clk;                                        // pll_0_50:outclk_0 -> [in_fifo_used:clk, in_port_data:clk, in_port_dig_error:clk, in_port_ec_flags:clk, in_port_freq_cnt:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_50_outclk0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, out_port_batnum:clk, out_port_ctrl:clk, out_port_lut_adr:clk, out_port_lut_data:clk, out_port_prodnum:clk, product_info_0:clk, rst_controller:clk, rst_controller_001:clk, sysid_qsys_0:clock, timer_0:clk, uart_0:clk]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001:reset_in1]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [19:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [19:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_product_info_0_avalon_slave_0_chipselect;  // mm_interconnect_0:product_info_0_avalon_slave_0_chipselect -> product_info_0:chipselect_n
	wire  [31:0] mm_interconnect_0_product_info_0_avalon_slave_0_readdata;    // product_info_0:av_data_read -> mm_interconnect_0:product_info_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_product_info_0_avalon_slave_0_address;     // mm_interconnect_0:product_info_0_avalon_slave_0_address -> product_info_0:av_address
	wire         mm_interconnect_0_product_info_0_avalon_slave_0_read;        // mm_interconnect_0:product_info_0_avalon_slave_0_read -> product_info_0:read_n
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_in_fifo_used_s1_readdata;                  // in_fifo_used:readdata -> mm_interconnect_0:in_fifo_used_s1_readdata
	wire   [1:0] mm_interconnect_0_in_fifo_used_s1_address;                   // mm_interconnect_0:in_fifo_used_s1_address -> in_fifo_used:address
	wire  [31:0] mm_interconnect_0_in_port_data_s1_readdata;                  // in_port_data:readdata -> mm_interconnect_0:in_port_data_s1_readdata
	wire   [1:0] mm_interconnect_0_in_port_data_s1_address;                   // mm_interconnect_0:in_port_data_s1_address -> in_port_data:address
	wire  [31:0] mm_interconnect_0_in_port_ec_flags_s1_readdata;              // in_port_ec_flags:readdata -> mm_interconnect_0:in_port_ec_flags_s1_readdata
	wire   [1:0] mm_interconnect_0_in_port_ec_flags_s1_address;               // mm_interconnect_0:in_port_ec_flags_s1_address -> in_port_ec_flags:address
	wire         mm_interconnect_0_out_port_ctrl_s1_chipselect;               // mm_interconnect_0:out_port_ctrl_s1_chipselect -> out_port_ctrl:chipselect
	wire  [31:0] mm_interconnect_0_out_port_ctrl_s1_readdata;                 // out_port_ctrl:readdata -> mm_interconnect_0:out_port_ctrl_s1_readdata
	wire   [1:0] mm_interconnect_0_out_port_ctrl_s1_address;                  // mm_interconnect_0:out_port_ctrl_s1_address -> out_port_ctrl:address
	wire         mm_interconnect_0_out_port_ctrl_s1_write;                    // mm_interconnect_0:out_port_ctrl_s1_write -> out_port_ctrl:write_n
	wire  [31:0] mm_interconnect_0_out_port_ctrl_s1_writedata;                // mm_interconnect_0:out_port_ctrl_s1_writedata -> out_port_ctrl:writedata
	wire  [31:0] mm_interconnect_0_in_port_dig_error_s1_readdata;             // in_port_dig_error:readdata -> mm_interconnect_0:in_port_dig_error_s1_readdata
	wire   [1:0] mm_interconnect_0_in_port_dig_error_s1_address;              // mm_interconnect_0:in_port_dig_error_s1_address -> in_port_dig_error:address
	wire         mm_interconnect_0_uart_0_s1_chipselect;                      // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                        // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                         // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                            // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                   // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                           // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                       // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_out_port_prodnum_s1_chipselect;            // mm_interconnect_0:out_port_prodnum_s1_chipselect -> out_port_prodnum:chipselect
	wire  [31:0] mm_interconnect_0_out_port_prodnum_s1_readdata;              // out_port_prodnum:readdata -> mm_interconnect_0:out_port_prodnum_s1_readdata
	wire   [1:0] mm_interconnect_0_out_port_prodnum_s1_address;               // mm_interconnect_0:out_port_prodnum_s1_address -> out_port_prodnum:address
	wire         mm_interconnect_0_out_port_prodnum_s1_write;                 // mm_interconnect_0:out_port_prodnum_s1_write -> out_port_prodnum:write_n
	wire  [31:0] mm_interconnect_0_out_port_prodnum_s1_writedata;             // mm_interconnect_0:out_port_prodnum_s1_writedata -> out_port_prodnum:writedata
	wire         mm_interconnect_0_out_port_batnum_s1_chipselect;             // mm_interconnect_0:out_port_batnum_s1_chipselect -> out_port_batnum:chipselect
	wire  [31:0] mm_interconnect_0_out_port_batnum_s1_readdata;               // out_port_batnum:readdata -> mm_interconnect_0:out_port_batnum_s1_readdata
	wire   [1:0] mm_interconnect_0_out_port_batnum_s1_address;                // mm_interconnect_0:out_port_batnum_s1_address -> out_port_batnum:address
	wire         mm_interconnect_0_out_port_batnum_s1_write;                  // mm_interconnect_0:out_port_batnum_s1_write -> out_port_batnum:write_n
	wire  [31:0] mm_interconnect_0_out_port_batnum_s1_writedata;              // mm_interconnect_0:out_port_batnum_s1_writedata -> out_port_batnum:writedata
	wire         mm_interconnect_0_out_port_lut_data_s1_chipselect;           // mm_interconnect_0:out_port_lut_data_s1_chipselect -> out_port_lut_data:chipselect
	wire  [31:0] mm_interconnect_0_out_port_lut_data_s1_readdata;             // out_port_lut_data:readdata -> mm_interconnect_0:out_port_lut_data_s1_readdata
	wire   [1:0] mm_interconnect_0_out_port_lut_data_s1_address;              // mm_interconnect_0:out_port_lut_data_s1_address -> out_port_lut_data:address
	wire         mm_interconnect_0_out_port_lut_data_s1_write;                // mm_interconnect_0:out_port_lut_data_s1_write -> out_port_lut_data:write_n
	wire  [31:0] mm_interconnect_0_out_port_lut_data_s1_writedata;            // mm_interconnect_0:out_port_lut_data_s1_writedata -> out_port_lut_data:writedata
	wire         mm_interconnect_0_out_port_lut_adr_s1_chipselect;            // mm_interconnect_0:out_port_lut_adr_s1_chipselect -> out_port_lut_adr:chipselect
	wire  [31:0] mm_interconnect_0_out_port_lut_adr_s1_readdata;              // out_port_lut_adr:readdata -> mm_interconnect_0:out_port_lut_adr_s1_readdata
	wire   [1:0] mm_interconnect_0_out_port_lut_adr_s1_address;               // mm_interconnect_0:out_port_lut_adr_s1_address -> out_port_lut_adr:address
	wire         mm_interconnect_0_out_port_lut_adr_s1_write;                 // mm_interconnect_0:out_port_lut_adr_s1_write -> out_port_lut_adr:write_n
	wire  [31:0] mm_interconnect_0_out_port_lut_adr_s1_writedata;             // mm_interconnect_0:out_port_lut_adr_s1_writedata -> out_port_lut_adr:writedata
	wire  [31:0] mm_interconnect_0_in_port_freq_cnt_s1_readdata;              // in_port_freq_cnt:readdata -> mm_interconnect_0:in_port_freq_cnt_s1_readdata
	wire   [1:0] mm_interconnect_0_in_port_freq_cnt_s1_address;               // mm_interconnect_0:in_port_freq_cnt_s1_address -> in_port_freq_cnt:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // uart_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [in_fifo_used:reset_n, in_port_data:reset_n, in_port_dig_error:reset_n, in_port_ec_flags:reset_n, in_port_freq_cnt:reset_n, mm_interconnect_0:product_info_0_clock_reset_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, out_port_batnum:reset_n, out_port_ctrl:reset_n, out_port_lut_adr:reset_n, out_port_lut_data:reset_n, out_port_prodnum:reset_n, product_info_0:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n, timer_0:reset_n, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]

	q_sys_in_fifo_used in_fifo_used (
		.clk      (pll_0_50_outclk0_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_in_fifo_used_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_fifo_used_s1_readdata), //                    .readdata
		.in_port  (in_fifo_used_external_connection_export)     // external_connection.export
	);

	q_sys_in_port_data in_port_data (
		.clk      (pll_0_50_outclk0_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_in_port_data_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_port_data_s1_readdata), //                    .readdata
		.in_port  (in_port_data_external_connection_export)     // external_connection.export
	);

	q_sys_in_port_dig_error in_port_dig_error (
		.clk      (pll_0_50_outclk0_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_in_port_dig_error_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_port_dig_error_s1_readdata), //                    .readdata
		.in_port  (in_port_dig_error_external_connection_export)     // external_connection.export
	);

	q_sys_in_port_ec_flags in_port_ec_flags (
		.clk      (pll_0_50_outclk0_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_in_port_ec_flags_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_port_ec_flags_s1_readdata), //                    .readdata
		.in_port  (in_port_ec_flags_external_connection_export)     // external_connection.export
	);

	q_sys_in_port_freq_cnt in_port_freq_cnt (
		.clk      (pll_0_50_outclk0_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_in_port_freq_cnt_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_in_port_freq_cnt_s1_readdata), //                    .readdata
		.in_port  (in_port_freq_cnt_external_connection_export)     // external_connection.export
	);

	q_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_0_50_outclk0_clk),                                        //               clk.clk
		.rst_n          (~nios2_gen2_0_debug_reset_request_reset),                     //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	q_sys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_0_50_outclk0_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	q_sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_0_50_outclk0_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	q_sys_out_port_batnum out_port_batnum (
		.clk        (pll_0_50_outclk0_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_out_port_batnum_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_port_batnum_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_port_batnum_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_port_batnum_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_port_batnum_s1_readdata),   //                    .readdata
		.out_port   (out_port_batnum_external_connection_export)       // external_connection.export
	);

	q_sys_out_port_ctrl out_port_ctrl (
		.clk        (pll_0_50_outclk0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_out_port_ctrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_port_ctrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_port_ctrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_port_ctrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_port_ctrl_s1_readdata),   //                    .readdata
		.out_port   (out_port_ctrl_external_connection_export)       // external_connection.export
	);

	q_sys_out_port_lut_adr out_port_lut_adr (
		.clk        (pll_0_50_outclk0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_out_port_lut_adr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_port_lut_adr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_port_lut_adr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_port_lut_adr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_port_lut_adr_s1_readdata),   //                    .readdata
		.out_port   (out_port_lut_adr_external_connection_export)       // external_connection.export
	);

	q_sys_out_port_lut_data out_port_lut_data (
		.clk        (pll_0_50_outclk0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_out_port_lut_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_port_lut_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_port_lut_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_port_lut_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_port_lut_data_s1_readdata),   //                    .readdata
		.out_port   (out_port_lut_data_external_connection_export)       // external_connection.export
	);

	q_sys_out_port_batnum out_port_prodnum (
		.clk        (pll_0_50_outclk0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_out_port_prodnum_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_out_port_prodnum_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_out_port_prodnum_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_out_port_prodnum_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_out_port_prodnum_s1_readdata),   //                    .readdata
		.out_port   (out_port_prodnum_external_connection_export)       // external_connection.export
	);

	q_sys_pll_0_50 pll_0_50 (
		.refclk   (clk_clk),              //  refclk.clk
		.rst      (~reset_reset_n),       //   reset.reset
		.outclk_0 (pll_0_50_outclk0_clk), // outclk0.clk
		.locked   ()                      // (terminated)
	);

	product_info product_info_0 (
		.clk          (pll_0_50_outclk0_clk),                                        //       clock_reset.clk
		.reset_n      (~rst_controller_reset_out_reset),                             // clock_reset_reset.reset_n
		.chipselect_n (~mm_interconnect_0_product_info_0_avalon_slave_0_chipselect), //    avalon_slave_0.chipselect_n
		.read_n       (~mm_interconnect_0_product_info_0_avalon_slave_0_read),       //                  .read_n
		.av_data_read (mm_interconnect_0_product_info_0_avalon_slave_0_readdata),    //                  .readdata
		.av_address   (mm_interconnect_0_product_info_0_avalon_slave_0_address)      //                  .address
	);

	q_sys_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_0_50_outclk0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	q_sys_timer_0 timer_0 (
		.clk        (pll_0_50_outclk0_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	q_sys_uart_0 uart_0 (
		.clk           (pll_0_50_outclk0_clk),                      //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	q_sys_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_50_outclk0_clk                                         (pll_0_50_outclk0_clk),                                        //                                       pll_0_50_outclk0.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset                (nios2_gen2_0_debug_reset_request_reset),                      //                jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                          //               nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.product_info_0_clock_reset_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // product_info_0_clock_reset_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                             (nios2_gen2_0_data_master_address),                            //                               nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                         (nios2_gen2_0_data_master_waitrequest),                        //                                                       .waitrequest
		.nios2_gen2_0_data_master_byteenable                          (nios2_gen2_0_data_master_byteenable),                         //                                                       .byteenable
		.nios2_gen2_0_data_master_read                                (nios2_gen2_0_data_master_read),                               //                                                       .read
		.nios2_gen2_0_data_master_readdata                            (nios2_gen2_0_data_master_readdata),                           //                                                       .readdata
		.nios2_gen2_0_data_master_write                               (nios2_gen2_0_data_master_write),                              //                                                       .write
		.nios2_gen2_0_data_master_writedata                           (nios2_gen2_0_data_master_writedata),                          //                                                       .writedata
		.nios2_gen2_0_data_master_debugaccess                         (nios2_gen2_0_data_master_debugaccess),                        //                                                       .debugaccess
		.nios2_gen2_0_instruction_master_address                      (nios2_gen2_0_instruction_master_address),                     //                        nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                  (nios2_gen2_0_instruction_master_waitrequest),                 //                                                       .waitrequest
		.nios2_gen2_0_instruction_master_read                         (nios2_gen2_0_instruction_master_read),                        //                                                       .read
		.nios2_gen2_0_instruction_master_readdata                     (nios2_gen2_0_instruction_master_readdata),                    //                                                       .readdata
		.in_fifo_used_s1_address                                      (mm_interconnect_0_in_fifo_used_s1_address),                   //                                        in_fifo_used_s1.address
		.in_fifo_used_s1_readdata                                     (mm_interconnect_0_in_fifo_used_s1_readdata),                  //                                                       .readdata
		.in_port_data_s1_address                                      (mm_interconnect_0_in_port_data_s1_address),                   //                                        in_port_data_s1.address
		.in_port_data_s1_readdata                                     (mm_interconnect_0_in_port_data_s1_readdata),                  //                                                       .readdata
		.in_port_dig_error_s1_address                                 (mm_interconnect_0_in_port_dig_error_s1_address),              //                                   in_port_dig_error_s1.address
		.in_port_dig_error_s1_readdata                                (mm_interconnect_0_in_port_dig_error_s1_readdata),             //                                                       .readdata
		.in_port_ec_flags_s1_address                                  (mm_interconnect_0_in_port_ec_flags_s1_address),               //                                    in_port_ec_flags_s1.address
		.in_port_ec_flags_s1_readdata                                 (mm_interconnect_0_in_port_ec_flags_s1_readdata),              //                                                       .readdata
		.in_port_freq_cnt_s1_address                                  (mm_interconnect_0_in_port_freq_cnt_s1_address),               //                                    in_port_freq_cnt_s1.address
		.in_port_freq_cnt_s1_readdata                                 (mm_interconnect_0_in_port_freq_cnt_s1_readdata),              //                                                       .readdata
		.jtag_uart_0_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                          jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                       .write
		.jtag_uart_0_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                       .read
		.jtag_uart_0_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                       .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                       .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                       .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                       .chipselect
		.nios2_gen2_0_debug_mem_slave_address                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                           nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                                       .write
		.nios2_gen2_0_debug_mem_slave_read                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                                       .read
		.nios2_gen2_0_debug_mem_slave_readdata                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                                       .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                                       .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                                       .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                                       .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                                       .debugaccess
		.onchip_memory2_0_s1_address                                  (mm_interconnect_0_onchip_memory2_0_s1_address),               //                                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                    (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                                       .write
		.onchip_memory2_0_s1_readdata                                 (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                                       .readdata
		.onchip_memory2_0_s1_writedata                                (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                                       .writedata
		.onchip_memory2_0_s1_byteenable                               (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                                       .byteenable
		.onchip_memory2_0_s1_chipselect                               (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                                       .chipselect
		.onchip_memory2_0_s1_clken                                    (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                                       .clken
		.out_port_batnum_s1_address                                   (mm_interconnect_0_out_port_batnum_s1_address),                //                                     out_port_batnum_s1.address
		.out_port_batnum_s1_write                                     (mm_interconnect_0_out_port_batnum_s1_write),                  //                                                       .write
		.out_port_batnum_s1_readdata                                  (mm_interconnect_0_out_port_batnum_s1_readdata),               //                                                       .readdata
		.out_port_batnum_s1_writedata                                 (mm_interconnect_0_out_port_batnum_s1_writedata),              //                                                       .writedata
		.out_port_batnum_s1_chipselect                                (mm_interconnect_0_out_port_batnum_s1_chipselect),             //                                                       .chipselect
		.out_port_ctrl_s1_address                                     (mm_interconnect_0_out_port_ctrl_s1_address),                  //                                       out_port_ctrl_s1.address
		.out_port_ctrl_s1_write                                       (mm_interconnect_0_out_port_ctrl_s1_write),                    //                                                       .write
		.out_port_ctrl_s1_readdata                                    (mm_interconnect_0_out_port_ctrl_s1_readdata),                 //                                                       .readdata
		.out_port_ctrl_s1_writedata                                   (mm_interconnect_0_out_port_ctrl_s1_writedata),                //                                                       .writedata
		.out_port_ctrl_s1_chipselect                                  (mm_interconnect_0_out_port_ctrl_s1_chipselect),               //                                                       .chipselect
		.out_port_lut_adr_s1_address                                  (mm_interconnect_0_out_port_lut_adr_s1_address),               //                                    out_port_lut_adr_s1.address
		.out_port_lut_adr_s1_write                                    (mm_interconnect_0_out_port_lut_adr_s1_write),                 //                                                       .write
		.out_port_lut_adr_s1_readdata                                 (mm_interconnect_0_out_port_lut_adr_s1_readdata),              //                                                       .readdata
		.out_port_lut_adr_s1_writedata                                (mm_interconnect_0_out_port_lut_adr_s1_writedata),             //                                                       .writedata
		.out_port_lut_adr_s1_chipselect                               (mm_interconnect_0_out_port_lut_adr_s1_chipselect),            //                                                       .chipselect
		.out_port_lut_data_s1_address                                 (mm_interconnect_0_out_port_lut_data_s1_address),              //                                   out_port_lut_data_s1.address
		.out_port_lut_data_s1_write                                   (mm_interconnect_0_out_port_lut_data_s1_write),                //                                                       .write
		.out_port_lut_data_s1_readdata                                (mm_interconnect_0_out_port_lut_data_s1_readdata),             //                                                       .readdata
		.out_port_lut_data_s1_writedata                               (mm_interconnect_0_out_port_lut_data_s1_writedata),            //                                                       .writedata
		.out_port_lut_data_s1_chipselect                              (mm_interconnect_0_out_port_lut_data_s1_chipselect),           //                                                       .chipselect
		.out_port_prodnum_s1_address                                  (mm_interconnect_0_out_port_prodnum_s1_address),               //                                    out_port_prodnum_s1.address
		.out_port_prodnum_s1_write                                    (mm_interconnect_0_out_port_prodnum_s1_write),                 //                                                       .write
		.out_port_prodnum_s1_readdata                                 (mm_interconnect_0_out_port_prodnum_s1_readdata),              //                                                       .readdata
		.out_port_prodnum_s1_writedata                                (mm_interconnect_0_out_port_prodnum_s1_writedata),             //                                                       .writedata
		.out_port_prodnum_s1_chipselect                               (mm_interconnect_0_out_port_prodnum_s1_chipselect),            //                                                       .chipselect
		.product_info_0_avalon_slave_0_address                        (mm_interconnect_0_product_info_0_avalon_slave_0_address),     //                          product_info_0_avalon_slave_0.address
		.product_info_0_avalon_slave_0_read                           (mm_interconnect_0_product_info_0_avalon_slave_0_read),        //                                                       .read
		.product_info_0_avalon_slave_0_readdata                       (mm_interconnect_0_product_info_0_avalon_slave_0_readdata),    //                                                       .readdata
		.product_info_0_avalon_slave_0_chipselect                     (mm_interconnect_0_product_info_0_avalon_slave_0_chipselect),  //                                                       .chipselect
		.sysid_qsys_0_control_slave_address                           (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //                             sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                          (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                                       .readdata
		.timer_0_s1_address                                           (mm_interconnect_0_timer_0_s1_address),                        //                                             timer_0_s1.address
		.timer_0_s1_write                                             (mm_interconnect_0_timer_0_s1_write),                          //                                                       .write
		.timer_0_s1_readdata                                          (mm_interconnect_0_timer_0_s1_readdata),                       //                                                       .readdata
		.timer_0_s1_writedata                                         (mm_interconnect_0_timer_0_s1_writedata),                      //                                                       .writedata
		.timer_0_s1_chipselect                                        (mm_interconnect_0_timer_0_s1_chipselect),                     //                                                       .chipselect
		.uart_0_s1_address                                            (mm_interconnect_0_uart_0_s1_address),                         //                                              uart_0_s1.address
		.uart_0_s1_write                                              (mm_interconnect_0_uart_0_s1_write),                           //                                                       .write
		.uart_0_s1_read                                               (mm_interconnect_0_uart_0_s1_read),                            //                                                       .read
		.uart_0_s1_readdata                                           (mm_interconnect_0_uart_0_s1_readdata),                        //                                                       .readdata
		.uart_0_s1_writedata                                          (mm_interconnect_0_uart_0_s1_writedata),                       //                                                       .writedata
		.uart_0_s1_begintransfer                                      (mm_interconnect_0_uart_0_s1_begintransfer),                   //                                                       .begintransfer
		.uart_0_s1_chipselect                                         (mm_interconnect_0_uart_0_s1_chipselect)                       //                                                       .chipselect
	);

	q_sys_irq_mapper irq_mapper (
		.clk           (pll_0_50_outclk0_clk),               //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_50_outclk0_clk),               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_0_50_outclk0_clk),                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule

// q_sys_mSGDMA_0.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module q_sys_mSGDMA_0 (
		output wire         mm_bridge_slv_waitrequest,       //            mm_bridge_slv.waitrequest
		output wire [31:0]  mm_bridge_slv_readdata,          //                         .readdata
		output wire         mm_bridge_slv_readdatavalid,     //                         .readdatavalid
		input  wire [0:0]   mm_bridge_slv_burstcount,        //                         .burstcount
		input  wire [31:0]  mm_bridge_slv_writedata,         //                         .writedata
		input  wire [19:0]  mm_bridge_slv_address,           //                         .address
		input  wire         mm_bridge_slv_write,             //                         .write
		input  wire         mm_bridge_slv_read,              //                         .read
		input  wire [3:0]   mm_bridge_slv_byteenable,        //                         .byteenable
		input  wire         mm_bridge_slv_debugaccess,       //                         .debugaccess
		input  wire         reset_reset_n,                   //                    reset.reset_n
		input  wire         clk_clk,                         //                      clk.clk
		output wire [27:0]  dma_read_master_address,         //          dma_read_master.address
		output wire         dma_read_master_read,            //                         .read
		output wire [31:0]  dma_read_master_byteenable,      //                         .byteenable
		input  wire [255:0] dma_read_master_readdata,        //                         .readdata
		input  wire         dma_read_master_waitrequest,     //                         .waitrequest
		input  wire         dma_read_master_readdatavalid,   //                         .readdatavalid
		output wire [5:0]   dma_read_master_burstcount,      //                         .burstcount
		output wire [27:0]  dma_write_master_address,        //         dma_write_master.address
		output wire         dma_write_master_write,          //                         .write
		output wire [31:0]  dma_write_master_byteenable,     //                         .byteenable
		output wire [255:0] dma_write_master_writedata,      //                         .writedata
		input  wire         dma_write_master_waitrequest,    //                         .waitrequest
		output wire [5:0]   dma_write_master_burstcount,     //                         .burstcount
		output wire         dispatcher_write_csr_irq_irq,    // dispatcher_write_csr_irq.irq
		output wire         dispatcher_read_csr_irq_irq,     //  dispatcher_read_csr_irq.irq
		input  wire         clk_0_clk,                       //                    clk_0.clk
		input  wire         reset_0_reset_n,                 //                  reset_0.reset_n
		output wire         status_mon_out_cal_fail_mon,     //           status_mon_out.cal_fail_mon
		output wire         status_mon_out_cal_success_mon,  //                         .cal_success_mon
		output wire         status_mon_out_init_done_mon,    //                         .init_done_mon
		input  wire         status_mon_in_local_init_done,   //            status_mon_in.local_init_done
		input  wire         status_mon_in_local_cal_success, //                         .local_cal_success
		input  wire         status_mon_in_local_cal_fail,    //                         .local_cal_fail
		output wire         reset_source_reset_n             //             reset_source.reset_n
	);

	wire          prbs_pattern_generator_st_pattern_output_valid;                  // prbs_pattern_generator:src_valid -> timing_adapter:in_valid
	wire  [255:0] prbs_pattern_generator_st_pattern_output_data;                   // prbs_pattern_generator:src_data -> timing_adapter:in_data
	wire          prbs_pattern_generator_st_pattern_output_ready;                  // timing_adapter:in_ready -> prbs_pattern_generator:src_ready
	wire          timing_adapter_out_valid;                                        // timing_adapter:out_valid -> dma_write_master:snk_valid
	wire  [255:0] timing_adapter_out_data;                                         // timing_adapter:out_data -> dma_write_master:snk_data
	wire          timing_adapter_out_ready;                                        // dma_write_master:snk_ready -> timing_adapter:out_ready
	wire          dispatcher_write_write_command_source_valid;                     // dispatcher_write:src_write_master_valid -> dma_write_master:snk_command_valid
	wire  [255:0] dispatcher_write_write_command_source_data;                      // dispatcher_write:src_write_master_data -> dma_write_master:snk_command_data
	wire          dispatcher_write_write_command_source_ready;                     // dma_write_master:snk_command_ready -> dispatcher_write:src_write_master_ready
	wire          dma_write_master_response_source_valid;                          // dma_write_master:src_response_valid -> dispatcher_write:snk_write_master_valid
	wire  [255:0] dma_write_master_response_source_data;                           // dma_write_master:src_response_data -> dispatcher_write:snk_write_master_data
	wire          dma_write_master_response_source_ready;                          // dispatcher_write:snk_write_master_ready -> dma_write_master:src_response_ready
	wire          dma_read_master_data_source_valid;                               // dma_read_master:src_valid -> prbs_pattern_checker:snk_valid
	wire  [255:0] dma_read_master_data_source_data;                                // dma_read_master:src_data -> prbs_pattern_checker:snk_data
	wire          dma_read_master_data_source_ready;                               // prbs_pattern_checker:snk_ready -> dma_read_master:src_ready
	wire          dispatcher_read_read_command_source_valid;                       // dispatcher_read:src_read_master_valid -> dma_read_master:snk_command_valid
	wire  [255:0] dispatcher_read_read_command_source_data;                        // dispatcher_read:src_read_master_data -> dma_read_master:snk_command_data
	wire          dispatcher_read_read_command_source_ready;                       // dma_read_master:snk_command_ready -> dispatcher_read:src_read_master_ready
	wire          dma_read_master_response_source_valid;                           // dma_read_master:src_response_valid -> dispatcher_read:snk_read_master_valid
	wire  [255:0] dma_read_master_response_source_data;                            // dma_read_master:src_response_data -> dispatcher_read:snk_read_master_data
	wire          dma_read_master_response_source_ready;                           // dispatcher_read:snk_read_master_ready -> dma_read_master:src_response_ready
	wire          mm_bridge_slv_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_slv_m0_waitrequest -> mm_bridge_slv:m0_waitrequest
	wire   [31:0] mm_bridge_slv_m0_readdata;                                       // mm_interconnect_0:mm_bridge_slv_m0_readdata -> mm_bridge_slv:m0_readdata
	wire          mm_bridge_slv_m0_debugaccess;                                    // mm_bridge_slv:m0_debugaccess -> mm_interconnect_0:mm_bridge_slv_m0_debugaccess
	wire   [19:0] mm_bridge_slv_m0_address;                                        // mm_bridge_slv:m0_address -> mm_interconnect_0:mm_bridge_slv_m0_address
	wire          mm_bridge_slv_m0_read;                                           // mm_bridge_slv:m0_read -> mm_interconnect_0:mm_bridge_slv_m0_read
	wire    [3:0] mm_bridge_slv_m0_byteenable;                                     // mm_bridge_slv:m0_byteenable -> mm_interconnect_0:mm_bridge_slv_m0_byteenable
	wire          mm_bridge_slv_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_slv_m0_readdatavalid -> mm_bridge_slv:m0_readdatavalid
	wire   [31:0] mm_bridge_slv_m0_writedata;                                      // mm_bridge_slv:m0_writedata -> mm_interconnect_0:mm_bridge_slv_m0_writedata
	wire          mm_bridge_slv_m0_write;                                          // mm_bridge_slv:m0_write -> mm_interconnect_0:mm_bridge_slv_m0_write
	wire    [0:0] mm_bridge_slv_m0_burstcount;                                     // mm_bridge_slv:m0_burstcount -> mm_interconnect_0:mm_bridge_slv_m0_burstcount
	wire   [31:0] mm_interconnect_0_prbs_pattern_generator_csr_readdata;           // prbs_pattern_generator:csr_readdata -> mm_interconnect_0:prbs_pattern_generator_csr_readdata
	wire    [2:0] mm_interconnect_0_prbs_pattern_generator_csr_address;            // mm_interconnect_0:prbs_pattern_generator_csr_address -> prbs_pattern_generator:csr_address
	wire          mm_interconnect_0_prbs_pattern_generator_csr_read;               // mm_interconnect_0:prbs_pattern_generator_csr_read -> prbs_pattern_generator:csr_read
	wire    [3:0] mm_interconnect_0_prbs_pattern_generator_csr_byteenable;         // mm_interconnect_0:prbs_pattern_generator_csr_byteenable -> prbs_pattern_generator:csr_byteenable
	wire          mm_interconnect_0_prbs_pattern_generator_csr_write;              // mm_interconnect_0:prbs_pattern_generator_csr_write -> prbs_pattern_generator:csr_write
	wire   [31:0] mm_interconnect_0_prbs_pattern_generator_csr_writedata;          // mm_interconnect_0:prbs_pattern_generator_csr_writedata -> prbs_pattern_generator:csr_writedata
	wire   [31:0] mm_interconnect_0_dispatcher_write_csr_readdata;                 // dispatcher_write:csr_readdata -> mm_interconnect_0:dispatcher_write_CSR_readdata
	wire    [2:0] mm_interconnect_0_dispatcher_write_csr_address;                  // mm_interconnect_0:dispatcher_write_CSR_address -> dispatcher_write:csr_address
	wire          mm_interconnect_0_dispatcher_write_csr_read;                     // mm_interconnect_0:dispatcher_write_CSR_read -> dispatcher_write:csr_read
	wire    [3:0] mm_interconnect_0_dispatcher_write_csr_byteenable;               // mm_interconnect_0:dispatcher_write_CSR_byteenable -> dispatcher_write:csr_byteenable
	wire          mm_interconnect_0_dispatcher_write_csr_write;                    // mm_interconnect_0:dispatcher_write_CSR_write -> dispatcher_write:csr_write
	wire   [31:0] mm_interconnect_0_dispatcher_write_csr_writedata;                // mm_interconnect_0:dispatcher_write_CSR_writedata -> dispatcher_write:csr_writedata
	wire          mm_interconnect_0_dispatcher_write_descriptor_slave_waitrequest; // dispatcher_write:descriptor_waitrequest -> mm_interconnect_0:dispatcher_write_Descriptor_Slave_waitrequest
	wire   [15:0] mm_interconnect_0_dispatcher_write_descriptor_slave_byteenable;  // mm_interconnect_0:dispatcher_write_Descriptor_Slave_byteenable -> dispatcher_write:descriptor_byteenable
	wire          mm_interconnect_0_dispatcher_write_descriptor_slave_write;       // mm_interconnect_0:dispatcher_write_Descriptor_Slave_write -> dispatcher_write:descriptor_write
	wire  [127:0] mm_interconnect_0_dispatcher_write_descriptor_slave_writedata;   // mm_interconnect_0:dispatcher_write_Descriptor_Slave_writedata -> dispatcher_write:descriptor_writedata
	wire   [31:0] mm_interconnect_0_prbs_pattern_checker_csr_readdata;             // prbs_pattern_checker:csr_readdata -> mm_interconnect_0:prbs_pattern_checker_csr_readdata
	wire    [3:0] mm_interconnect_0_prbs_pattern_checker_csr_address;              // mm_interconnect_0:prbs_pattern_checker_csr_address -> prbs_pattern_checker:csr_address
	wire          mm_interconnect_0_prbs_pattern_checker_csr_read;                 // mm_interconnect_0:prbs_pattern_checker_csr_read -> prbs_pattern_checker:csr_read
	wire    [3:0] mm_interconnect_0_prbs_pattern_checker_csr_byteenable;           // mm_interconnect_0:prbs_pattern_checker_csr_byteenable -> prbs_pattern_checker:csr_byteenable
	wire          mm_interconnect_0_prbs_pattern_checker_csr_write;                // mm_interconnect_0:prbs_pattern_checker_csr_write -> prbs_pattern_checker:csr_write
	wire   [31:0] mm_interconnect_0_prbs_pattern_checker_csr_writedata;            // mm_interconnect_0:prbs_pattern_checker_csr_writedata -> prbs_pattern_checker:csr_writedata
	wire   [31:0] mm_interconnect_0_dispatcher_read_csr_readdata;                  // dispatcher_read:csr_readdata -> mm_interconnect_0:dispatcher_read_CSR_readdata
	wire    [2:0] mm_interconnect_0_dispatcher_read_csr_address;                   // mm_interconnect_0:dispatcher_read_CSR_address -> dispatcher_read:csr_address
	wire          mm_interconnect_0_dispatcher_read_csr_read;                      // mm_interconnect_0:dispatcher_read_CSR_read -> dispatcher_read:csr_read
	wire    [3:0] mm_interconnect_0_dispatcher_read_csr_byteenable;                // mm_interconnect_0:dispatcher_read_CSR_byteenable -> dispatcher_read:csr_byteenable
	wire          mm_interconnect_0_dispatcher_read_csr_write;                     // mm_interconnect_0:dispatcher_read_CSR_write -> dispatcher_read:csr_write
	wire   [31:0] mm_interconnect_0_dispatcher_read_csr_writedata;                 // mm_interconnect_0:dispatcher_read_CSR_writedata -> dispatcher_read:csr_writedata
	wire          mm_interconnect_0_dispatcher_read_descriptor_slave_waitrequest;  // dispatcher_read:descriptor_waitrequest -> mm_interconnect_0:dispatcher_read_Descriptor_Slave_waitrequest
	wire   [15:0] mm_interconnect_0_dispatcher_read_descriptor_slave_byteenable;   // mm_interconnect_0:dispatcher_read_Descriptor_Slave_byteenable -> dispatcher_read:descriptor_byteenable
	wire          mm_interconnect_0_dispatcher_read_descriptor_slave_write;        // mm_interconnect_0:dispatcher_read_Descriptor_Slave_write -> dispatcher_read:descriptor_write
	wire  [127:0] mm_interconnect_0_dispatcher_read_descriptor_slave_writedata;    // mm_interconnect_0:dispatcher_read_Descriptor_Slave_writedata -> dispatcher_read:descriptor_writedata
	wire          mm_interconnect_0_status_mon_0_slv_chipselect;                   // mm_interconnect_0:status_mon_0_slv_chipselect -> status_mon_0:slv_cs_n
	wire   [31:0] mm_interconnect_0_status_mon_0_slv_readdata;                     // status_mon_0:slv_data_read -> mm_interconnect_0:status_mon_0_slv_readdata
	wire    [1:0] mm_interconnect_0_status_mon_0_slv_address;                      // mm_interconnect_0:status_mon_0_slv_address -> status_mon_0:slv_address
	wire          mm_interconnect_0_status_mon_0_slv_read;                         // mm_interconnect_0:status_mon_0_slv_read -> status_mon_0:slv_read_n
	wire          mm_interconnect_0_status_mon_0_slv_write;                        // mm_interconnect_0:status_mon_0_slv_write -> status_mon_0:slv_write_n
	wire   [31:0] mm_interconnect_0_status_mon_0_slv_writedata;                    // mm_interconnect_0:status_mon_0_slv_writedata -> status_mon_0:slv_data_write
	wire   [31:0] mm_interconnect_0_frequency_counter_0_csr_readdata;              // frequency_counter_0:csr_readdata -> mm_interconnect_0:frequency_counter_0_csr_readdata
	wire          mm_interconnect_0_frequency_counter_0_csr_waitrequest;           // frequency_counter_0:csr_waitrequest -> mm_interconnect_0:frequency_counter_0_csr_waitrequest
	wire    [3:0] mm_interconnect_0_frequency_counter_0_csr_address;               // mm_interconnect_0:frequency_counter_0_csr_address -> frequency_counter_0:csr_address
	wire          mm_interconnect_0_frequency_counter_0_csr_read;                  // mm_interconnect_0:frequency_counter_0_csr_read -> frequency_counter_0:csr_read
	wire          mm_interconnect_0_timer_0_s1_chipselect;                         // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire   [15:0] mm_interconnect_0_timer_0_s1_readdata;                           // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire    [2:0] mm_interconnect_0_timer_0_s1_address;                            // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire          mm_interconnect_0_timer_0_s1_write;                              // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire   [15:0] mm_interconnect_0_timer_0_s1_writedata;                          // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire          rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [dispatcher_read:reset, dispatcher_write:reset, dma_read_master:reset, dma_write_master:reset, mm_bridge_slv:reset, mm_interconnect_0:mm_bridge_slv_reset_reset_bridge_in_reset_reset, prbs_pattern_checker:reset, prbs_pattern_generator:reset, status_mon_0:slv_reset_n, timing_adapter:reset_n]
	wire          rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [frequency_counter_0:reset_n, mm_interconnect_0:frequency_counter_0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> frequency_counter_0:sample_reset_n
	wire          rst_controller_003_reset_out_reset;                              // rst_controller_003:reset_out -> [mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, timer_0:reset_n]

	mtm_prbs_pattern_generator #(
		.DATA_WIDTH (256),
		.PRBS_WIDTH (32)
	) prbs_pattern_generator (
		.clk            (clk_clk),                                                 //             clock.clk
		.reset          (rst_controller_reset_out_reset),                          //             reset.reset
		.csr_address    (mm_interconnect_0_prbs_pattern_generator_csr_address),    //               csr.address
		.csr_writedata  (mm_interconnect_0_prbs_pattern_generator_csr_writedata),  //                  .writedata
		.csr_write      (mm_interconnect_0_prbs_pattern_generator_csr_write),      //                  .write
		.csr_readdata   (mm_interconnect_0_prbs_pattern_generator_csr_readdata),   //                  .readdata
		.csr_read       (mm_interconnect_0_prbs_pattern_generator_csr_read),       //                  .read
		.csr_byteenable (mm_interconnect_0_prbs_pattern_generator_csr_byteenable), //                  .byteenable
		.src_data       (prbs_pattern_generator_st_pattern_output_data),           // st_pattern_output.data
		.src_valid      (prbs_pattern_generator_st_pattern_output_valid),          //                  .valid
		.src_ready      (prbs_pattern_generator_st_pattern_output_ready)           //                  .ready
	);

	mtm_prbs_pattern_checker #(
		.DATA_WIDTH (256),
		.PRBS_WIDTH (32)
	) prbs_pattern_checker (
		.clk            (clk_clk),                                               //            clock.clk
		.reset          (rst_controller_reset_out_reset),                        //            reset.reset
		.csr_address    (mm_interconnect_0_prbs_pattern_checker_csr_address),    //              csr.address
		.csr_writedata  (mm_interconnect_0_prbs_pattern_checker_csr_writedata),  //                 .writedata
		.csr_write      (mm_interconnect_0_prbs_pattern_checker_csr_write),      //                 .write
		.csr_readdata   (mm_interconnect_0_prbs_pattern_checker_csr_readdata),   //                 .readdata
		.csr_read       (mm_interconnect_0_prbs_pattern_checker_csr_read),       //                 .read
		.csr_byteenable (mm_interconnect_0_prbs_pattern_checker_csr_byteenable), //                 .byteenable
		.snk_data       (dma_read_master_data_source_data),                      // st_pattern_input.data
		.snk_valid      (dma_read_master_data_source_valid),                     //                 .valid
		.snk_ready      (dma_read_master_data_source_ready)                      //                 .ready
	);

	write_master #(
		.DATA_WIDTH                     (256),
		.LENGTH_WIDTH                   (31),
		.FIFO_DEPTH                     (128),
		.STRIDE_ENABLE                  (0),
		.BURST_ENABLE                   (1),
		.PACKET_ENABLE                  (0),
		.ERROR_ENABLE                   (0),
		.ERROR_WIDTH                    (8),
		.BYTE_ENABLE_WIDTH              (32),
		.BYTE_ENABLE_WIDTH_LOG2         (5),
		.ADDRESS_WIDTH                  (28),
		.FIFO_DEPTH_LOG2                (7),
		.SYMBOL_WIDTH                   (8),
		.NUMBER_OF_SYMBOLS              (32),
		.NUMBER_OF_SYMBOLS_LOG2         (5),
		.MAX_BURST_COUNT_WIDTH          (6),
		.UNALIGNED_ACCESSES_ENABLE      (0),
		.ONLY_FULL_ACCESS_ENABLE        (1),
		.BURST_WRAPPING_SUPPORT         (0),
		.PROGRAMMABLE_BURST_ENABLE      (0),
		.MAX_BURST_COUNT                (32),
		.FIFO_SPEED_OPTIMIZATION        (1),
		.STRIDE_WIDTH                   (1),
		.ACTUAL_BYTES_TRANSFERRED_WIDTH (32)
	) dma_write_master (
		.clk                (clk_clk),                                     //             Clock.clk
		.reset              (rst_controller_reset_out_reset),              //       Clock_reset.reset
		.master_address     (dma_write_master_address),                    // Data_Write_Master.address
		.master_write       (dma_write_master_write),                      //                  .write
		.master_byteenable  (dma_write_master_byteenable),                 //                  .byteenable
		.master_writedata   (dma_write_master_writedata),                  //                  .writedata
		.master_waitrequest (dma_write_master_waitrequest),                //                  .waitrequest
		.master_burstcount  (dma_write_master_burstcount),                 //                  .burstcount
		.snk_data           (timing_adapter_out_data),                     //         Data_Sink.data
		.snk_valid          (timing_adapter_out_valid),                    //                  .valid
		.snk_ready          (timing_adapter_out_ready),                    //                  .ready
		.snk_command_data   (dispatcher_write_write_command_source_data),  //      Command_Sink.data
		.snk_command_valid  (dispatcher_write_write_command_source_valid), //                  .valid
		.snk_command_ready  (dispatcher_write_write_command_source_ready), //                  .ready
		.src_response_data  (dma_write_master_response_source_data),       //   Response_Source.data
		.src_response_valid (dma_write_master_response_source_valid),      //                  .valid
		.src_response_ready (dma_write_master_response_source_ready),      //                  .ready
		.snk_sop            (1'b0),                                        //       (terminated)
		.snk_eop            (1'b0),                                        //       (terminated)
		.snk_empty          (5'b00000),                                    //       (terminated)
		.snk_error          (8'b00000000)                                  //       (terminated)
	);

	dispatcher #(
		.MODE                        (2),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_FIFO_DEPTH       (8),
		.ENHANCED_FEATURES           (0),
		.DESCRIPTOR_WIDTH            (128),
		.DESCRIPTOR_BYTEENABLE_WIDTH (16),
		.CSR_ADDRESS_WIDTH           (3)
	) dispatcher_write (
		.clk                     (clk_clk),                                                                                                                                                                                                                                                               //                clock.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                                                                                                                                                        //          clock_reset.reset
		.csr_writedata           (mm_interconnect_0_dispatcher_write_csr_writedata),                                                                                                                                                                                                                      //                  CSR.writedata
		.csr_write               (mm_interconnect_0_dispatcher_write_csr_write),                                                                                                                                                                                                                          //                     .write
		.csr_byteenable          (mm_interconnect_0_dispatcher_write_csr_byteenable),                                                                                                                                                                                                                     //                     .byteenable
		.csr_readdata            (mm_interconnect_0_dispatcher_write_csr_readdata),                                                                                                                                                                                                                       //                     .readdata
		.csr_read                (mm_interconnect_0_dispatcher_write_csr_read),                                                                                                                                                                                                                           //                     .read
		.csr_address             (mm_interconnect_0_dispatcher_write_csr_address),                                                                                                                                                                                                                        //                     .address
		.descriptor_write        (mm_interconnect_0_dispatcher_write_descriptor_slave_write),                                                                                                                                                                                                             //     Descriptor_Slave.write
		.descriptor_waitrequest  (mm_interconnect_0_dispatcher_write_descriptor_slave_waitrequest),                                                                                                                                                                                                       //                     .waitrequest
		.descriptor_writedata    (mm_interconnect_0_dispatcher_write_descriptor_slave_writedata),                                                                                                                                                                                                         //                     .writedata
		.descriptor_byteenable   (mm_interconnect_0_dispatcher_write_descriptor_slave_byteenable),                                                                                                                                                                                                        //                     .byteenable
		.src_write_master_data   (dispatcher_write_write_command_source_data),                                                                                                                                                                                                                            // Write_Command_Source.data
		.src_write_master_valid  (dispatcher_write_write_command_source_valid),                                                                                                                                                                                                                           //                     .valid
		.src_write_master_ready  (dispatcher_write_write_command_source_ready),                                                                                                                                                                                                                           //                     .ready
		.snk_write_master_data   (dma_write_master_response_source_data),                                                                                                                                                                                                                                 //  Write_Response_Sink.data
		.snk_write_master_valid  (dma_write_master_response_source_valid),                                                                                                                                                                                                                                //                     .valid
		.snk_write_master_ready  (dma_write_master_response_source_ready),                                                                                                                                                                                                                                //                     .ready
		.csr_irq                 (dispatcher_write_csr_irq_irq),                                                                                                                                                                                                                                          //              csr_irq.irq
		.src_response_data       (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_response_valid      (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_response_ready      (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.mm_response_waitrequest (),                                                                                                                                                                                                                                                                      //          (terminated)
		.mm_response_byteenable  (4'b0000),                                                                                                                                                                                                                                                               //          (terminated)
		.mm_response_address     (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.mm_response_readdata    (),                                                                                                                                                                                                                                                                      //          (terminated)
		.mm_response_read        (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.src_read_master_data    (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_read_master_valid   (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_read_master_ready   (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.snk_read_master_data    (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //          (terminated)
		.snk_read_master_valid   (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.snk_read_master_ready   ()                                                                                                                                                                                                                                                                       //          (terminated)
	);

	read_master #(
		.DATA_WIDTH                (256),
		.LENGTH_WIDTH              (31),
		.FIFO_DEPTH                (128),
		.STRIDE_ENABLE             (0),
		.BURST_ENABLE              (1),
		.PACKET_ENABLE             (0),
		.ERROR_ENABLE              (0),
		.ERROR_WIDTH               (8),
		.CHANNEL_ENABLE            (0),
		.CHANNEL_WIDTH             (8),
		.BYTE_ENABLE_WIDTH         (32),
		.BYTE_ENABLE_WIDTH_LOG2    (5),
		.ADDRESS_WIDTH             (28),
		.FIFO_DEPTH_LOG2           (7),
		.SYMBOL_WIDTH              (8),
		.NUMBER_OF_SYMBOLS         (32),
		.NUMBER_OF_SYMBOLS_LOG2    (5),
		.MAX_BURST_COUNT_WIDTH     (6),
		.UNALIGNED_ACCESSES_ENABLE (0),
		.ONLY_FULL_ACCESS_ENABLE   (1),
		.BURST_WRAPPING_SUPPORT    (0),
		.PROGRAMMABLE_BURST_ENABLE (0),
		.MAX_BURST_COUNT           (32),
		.FIFO_SPEED_OPTIMIZATION   (1),
		.STRIDE_WIDTH              (1)
	) dma_read_master (
		.clk                  (clk_clk),                                   //            Clock.clk
		.reset                (rst_controller_reset_out_reset),            //      Clock_reset.reset
		.master_address       (dma_read_master_address),                   // Data_Read_Master.address
		.master_read          (dma_read_master_read),                      //                 .read
		.master_byteenable    (dma_read_master_byteenable),                //                 .byteenable
		.master_readdata      (dma_read_master_readdata),                  //                 .readdata
		.master_waitrequest   (dma_read_master_waitrequest),               //                 .waitrequest
		.master_readdatavalid (dma_read_master_readdatavalid),             //                 .readdatavalid
		.master_burstcount    (dma_read_master_burstcount),                //                 .burstcount
		.src_data             (dma_read_master_data_source_data),          //      Data_Source.data
		.src_valid            (dma_read_master_data_source_valid),         //                 .valid
		.src_ready            (dma_read_master_data_source_ready),         //                 .ready
		.snk_command_data     (dispatcher_read_read_command_source_data),  //     Command_Sink.data
		.snk_command_valid    (dispatcher_read_read_command_source_valid), //                 .valid
		.snk_command_ready    (dispatcher_read_read_command_source_ready), //                 .ready
		.src_response_data    (dma_read_master_response_source_data),      //  Response_Source.data
		.src_response_valid   (dma_read_master_response_source_valid),     //                 .valid
		.src_response_ready   (dma_read_master_response_source_ready),     //                 .ready
		.src_sop              (),                                          //      (terminated)
		.src_eop              (),                                          //      (terminated)
		.src_empty            (),                                          //      (terminated)
		.src_error            (),                                          //      (terminated)
		.src_channel          ()                                           //      (terminated)
	);

	dispatcher #(
		.MODE                        (1),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_FIFO_DEPTH       (8),
		.ENHANCED_FEATURES           (0),
		.DESCRIPTOR_WIDTH            (128),
		.DESCRIPTOR_BYTEENABLE_WIDTH (16),
		.CSR_ADDRESS_WIDTH           (3)
	) dispatcher_read (
		.clk                     (clk_clk),                                                                                                                                                                                                                                                               //               clock.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                                                                                                                                                        //         clock_reset.reset
		.csr_writedata           (mm_interconnect_0_dispatcher_read_csr_writedata),                                                                                                                                                                                                                       //                 CSR.writedata
		.csr_write               (mm_interconnect_0_dispatcher_read_csr_write),                                                                                                                                                                                                                           //                    .write
		.csr_byteenable          (mm_interconnect_0_dispatcher_read_csr_byteenable),                                                                                                                                                                                                                      //                    .byteenable
		.csr_readdata            (mm_interconnect_0_dispatcher_read_csr_readdata),                                                                                                                                                                                                                        //                    .readdata
		.csr_read                (mm_interconnect_0_dispatcher_read_csr_read),                                                                                                                                                                                                                            //                    .read
		.csr_address             (mm_interconnect_0_dispatcher_read_csr_address),                                                                                                                                                                                                                         //                    .address
		.descriptor_write        (mm_interconnect_0_dispatcher_read_descriptor_slave_write),                                                                                                                                                                                                              //    Descriptor_Slave.write
		.descriptor_waitrequest  (mm_interconnect_0_dispatcher_read_descriptor_slave_waitrequest),                                                                                                                                                                                                        //                    .waitrequest
		.descriptor_writedata    (mm_interconnect_0_dispatcher_read_descriptor_slave_writedata),                                                                                                                                                                                                          //                    .writedata
		.descriptor_byteenable   (mm_interconnect_0_dispatcher_read_descriptor_slave_byteenable),                                                                                                                                                                                                         //                    .byteenable
		.src_read_master_data    (dispatcher_read_read_command_source_data),                                                                                                                                                                                                                              // Read_Command_Source.data
		.src_read_master_valid   (dispatcher_read_read_command_source_valid),                                                                                                                                                                                                                             //                    .valid
		.src_read_master_ready   (dispatcher_read_read_command_source_ready),                                                                                                                                                                                                                             //                    .ready
		.snk_read_master_data    (dma_read_master_response_source_data),                                                                                                                                                                                                                                  //  Read_Response_Sink.data
		.snk_read_master_valid   (dma_read_master_response_source_valid),                                                                                                                                                                                                                                 //                    .valid
		.snk_read_master_ready   (dma_read_master_response_source_ready),                                                                                                                                                                                                                                 //                    .ready
		.csr_irq                 (dispatcher_read_csr_irq_irq),                                                                                                                                                                                                                                           //             csr_irq.irq
		.src_response_data       (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_response_valid      (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_response_ready      (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.mm_response_waitrequest (),                                                                                                                                                                                                                                                                      //         (terminated)
		.mm_response_byteenable  (4'b0000),                                                                                                                                                                                                                                                               //         (terminated)
		.mm_response_address     (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.mm_response_readdata    (),                                                                                                                                                                                                                                                                      //         (terminated)
		.mm_response_read        (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.src_write_master_data   (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_write_master_valid  (),                                                                                                                                                                                                                                                                      //         (terminated)
		.src_write_master_ready  (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.snk_write_master_data   (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.snk_write_master_valid  (1'b0),                                                                                                                                                                                                                                                                  //         (terminated)
		.snk_write_master_ready  ()                                                                                                                                                                                                                                                                       //         (terminated)
	);

	q_sys_mSGDMA_0_timing_adapter timing_adapter (
		.clk       (clk_clk),                                        //   clk.clk
		.reset_n   (~rst_controller_reset_out_reset),                // reset.reset_n
		.in_data   (prbs_pattern_generator_st_pattern_output_data),  //    in.data
		.in_valid  (prbs_pattern_generator_st_pattern_output_valid), //      .valid
		.in_ready  (prbs_pattern_generator_st_pattern_output_ready), //      .ready
		.out_data  (timing_adapter_out_data),                        //   out.data
		.out_valid (timing_adapter_out_valid),                       //      .valid
		.out_ready (timing_adapter_out_ready)                        //      .ready
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (20),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_slv (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (mm_bridge_slv_waitrequest),      //    s0.waitrequest
		.s0_readdata      (mm_bridge_slv_readdata),         //      .readdata
		.s0_readdatavalid (mm_bridge_slv_readdatavalid),    //      .readdatavalid
		.s0_burstcount    (mm_bridge_slv_burstcount),       //      .burstcount
		.s0_writedata     (mm_bridge_slv_writedata),        //      .writedata
		.s0_address       (mm_bridge_slv_address),          //      .address
		.s0_write         (mm_bridge_slv_write),            //      .write
		.s0_read          (mm_bridge_slv_read),             //      .read
		.s0_byteenable    (mm_bridge_slv_byteenable),       //      .byteenable
		.s0_debugaccess   (mm_bridge_slv_debugaccess),      //      .debugaccess
		.m0_waitrequest   (mm_bridge_slv_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_slv_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_slv_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_slv_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_slv_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_slv_m0_address),       //      .address
		.m0_write         (mm_bridge_slv_m0_write),         //      .write
		.m0_read          (mm_bridge_slv_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_slv_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_slv_m0_debugaccess),   //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	status_mon status_mon_0 (
		.slv_read_n        (~mm_interconnect_0_status_mon_0_slv_read),       //          slv.read_n
		.slv_write_n       (~mm_interconnect_0_status_mon_0_slv_write),      //             .write_n
		.slv_address       (mm_interconnect_0_status_mon_0_slv_address),     //             .address
		.slv_cs_n          (~mm_interconnect_0_status_mon_0_slv_chipselect), //             .chipselect_n
		.slv_data_write    (mm_interconnect_0_status_mon_0_slv_writedata),   //             .writedata
		.slv_data_read     (mm_interconnect_0_status_mon_0_slv_readdata),    //             .readdata
		.cal_fail_mon      (status_mon_out_cal_fail_mon),                    //  conduit_end.export
		.cal_success_mon   (status_mon_out_cal_success_mon),                 //             .export
		.init_done_mon     (status_mon_out_init_done_mon),                   //             .export
		.reset_out_n       (reset_source_reset_n),                           // reset_source.reset_n
		.slv_clk           (clk_clk),                                        //        clock.clk
		.slv_reset_n       (~rst_controller_reset_out_reset),                //      reset_n.reset_n
		.local_init_done   (status_mon_in_local_init_done),                  //       status.local_init_done
		.local_cal_success (status_mon_in_local_cal_success),                //             .local_cal_success
		.local_cal_fail    (status_mon_in_local_cal_fail)                    //             .local_cal_fail
	);

	frequency_counter #(
		.SYSTEM_CLK_FREQ_PICO_SEC (20000)
	) frequency_counter_0 (
		.reset_n         (~rst_controller_001_reset_out_reset),                   //          reset.reset_n
		.clk             (clk_0_clk),                                             //          clock.clk
		.csr_address     (mm_interconnect_0_frequency_counter_0_csr_address),     //            csr.address
		.csr_read        (mm_interconnect_0_frequency_counter_0_csr_read),        //               .read
		.csr_readdata    (mm_interconnect_0_frequency_counter_0_csr_readdata),    //               .readdata
		.csr_waitrequest (mm_interconnect_0_frequency_counter_0_csr_waitrequest), //               .waitrequest
		.sample_clk      (clk_clk),                                               //     sample_clk.clk
		.sample_reset_n  (~rst_controller_002_reset_out_reset)                    // sample_reset_n.reset_n
	);

	q_sys_mSGDMA_0_timer_0 timer_0 (
		.clk        (clk_0_clk),                               //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        ()                                         //   irq.irq
	);

	q_sys_mSGDMA_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                           (clk_clk),                                                         //                                         clk_clk.clk
		.clk_0_clk_clk                                         (clk_0_clk),                                                       //                                       clk_0_clk.clk
		.frequency_counter_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                              // frequency_counter_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_slv_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                  //       mm_bridge_slv_reset_reset_bridge_in_reset.reset
		.timer_0_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                              //             timer_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_slv_m0_address                              (mm_bridge_slv_m0_address),                                        //                                mm_bridge_slv_m0.address
		.mm_bridge_slv_m0_waitrequest                          (mm_bridge_slv_m0_waitrequest),                                    //                                                .waitrequest
		.mm_bridge_slv_m0_burstcount                           (mm_bridge_slv_m0_burstcount),                                     //                                                .burstcount
		.mm_bridge_slv_m0_byteenable                           (mm_bridge_slv_m0_byteenable),                                     //                                                .byteenable
		.mm_bridge_slv_m0_read                                 (mm_bridge_slv_m0_read),                                           //                                                .read
		.mm_bridge_slv_m0_readdata                             (mm_bridge_slv_m0_readdata),                                       //                                                .readdata
		.mm_bridge_slv_m0_readdatavalid                        (mm_bridge_slv_m0_readdatavalid),                                  //                                                .readdatavalid
		.mm_bridge_slv_m0_write                                (mm_bridge_slv_m0_write),                                          //                                                .write
		.mm_bridge_slv_m0_writedata                            (mm_bridge_slv_m0_writedata),                                      //                                                .writedata
		.mm_bridge_slv_m0_debugaccess                          (mm_bridge_slv_m0_debugaccess),                                    //                                                .debugaccess
		.dispatcher_read_CSR_address                           (mm_interconnect_0_dispatcher_read_csr_address),                   //                             dispatcher_read_CSR.address
		.dispatcher_read_CSR_write                             (mm_interconnect_0_dispatcher_read_csr_write),                     //                                                .write
		.dispatcher_read_CSR_read                              (mm_interconnect_0_dispatcher_read_csr_read),                      //                                                .read
		.dispatcher_read_CSR_readdata                          (mm_interconnect_0_dispatcher_read_csr_readdata),                  //                                                .readdata
		.dispatcher_read_CSR_writedata                         (mm_interconnect_0_dispatcher_read_csr_writedata),                 //                                                .writedata
		.dispatcher_read_CSR_byteenable                        (mm_interconnect_0_dispatcher_read_csr_byteenable),                //                                                .byteenable
		.dispatcher_read_Descriptor_Slave_write                (mm_interconnect_0_dispatcher_read_descriptor_slave_write),        //                dispatcher_read_Descriptor_Slave.write
		.dispatcher_read_Descriptor_Slave_writedata            (mm_interconnect_0_dispatcher_read_descriptor_slave_writedata),    //                                                .writedata
		.dispatcher_read_Descriptor_Slave_byteenable           (mm_interconnect_0_dispatcher_read_descriptor_slave_byteenable),   //                                                .byteenable
		.dispatcher_read_Descriptor_Slave_waitrequest          (mm_interconnect_0_dispatcher_read_descriptor_slave_waitrequest),  //                                                .waitrequest
		.dispatcher_write_CSR_address                          (mm_interconnect_0_dispatcher_write_csr_address),                  //                            dispatcher_write_CSR.address
		.dispatcher_write_CSR_write                            (mm_interconnect_0_dispatcher_write_csr_write),                    //                                                .write
		.dispatcher_write_CSR_read                             (mm_interconnect_0_dispatcher_write_csr_read),                     //                                                .read
		.dispatcher_write_CSR_readdata                         (mm_interconnect_0_dispatcher_write_csr_readdata),                 //                                                .readdata
		.dispatcher_write_CSR_writedata                        (mm_interconnect_0_dispatcher_write_csr_writedata),                //                                                .writedata
		.dispatcher_write_CSR_byteenable                       (mm_interconnect_0_dispatcher_write_csr_byteenable),               //                                                .byteenable
		.dispatcher_write_Descriptor_Slave_write               (mm_interconnect_0_dispatcher_write_descriptor_slave_write),       //               dispatcher_write_Descriptor_Slave.write
		.dispatcher_write_Descriptor_Slave_writedata           (mm_interconnect_0_dispatcher_write_descriptor_slave_writedata),   //                                                .writedata
		.dispatcher_write_Descriptor_Slave_byteenable          (mm_interconnect_0_dispatcher_write_descriptor_slave_byteenable),  //                                                .byteenable
		.dispatcher_write_Descriptor_Slave_waitrequest         (mm_interconnect_0_dispatcher_write_descriptor_slave_waitrequest), //                                                .waitrequest
		.frequency_counter_0_csr_address                       (mm_interconnect_0_frequency_counter_0_csr_address),               //                         frequency_counter_0_csr.address
		.frequency_counter_0_csr_read                          (mm_interconnect_0_frequency_counter_0_csr_read),                  //                                                .read
		.frequency_counter_0_csr_readdata                      (mm_interconnect_0_frequency_counter_0_csr_readdata),              //                                                .readdata
		.frequency_counter_0_csr_waitrequest                   (mm_interconnect_0_frequency_counter_0_csr_waitrequest),           //                                                .waitrequest
		.prbs_pattern_checker_csr_address                      (mm_interconnect_0_prbs_pattern_checker_csr_address),              //                        prbs_pattern_checker_csr.address
		.prbs_pattern_checker_csr_write                        (mm_interconnect_0_prbs_pattern_checker_csr_write),                //                                                .write
		.prbs_pattern_checker_csr_read                         (mm_interconnect_0_prbs_pattern_checker_csr_read),                 //                                                .read
		.prbs_pattern_checker_csr_readdata                     (mm_interconnect_0_prbs_pattern_checker_csr_readdata),             //                                                .readdata
		.prbs_pattern_checker_csr_writedata                    (mm_interconnect_0_prbs_pattern_checker_csr_writedata),            //                                                .writedata
		.prbs_pattern_checker_csr_byteenable                   (mm_interconnect_0_prbs_pattern_checker_csr_byteenable),           //                                                .byteenable
		.prbs_pattern_generator_csr_address                    (mm_interconnect_0_prbs_pattern_generator_csr_address),            //                      prbs_pattern_generator_csr.address
		.prbs_pattern_generator_csr_write                      (mm_interconnect_0_prbs_pattern_generator_csr_write),              //                                                .write
		.prbs_pattern_generator_csr_read                       (mm_interconnect_0_prbs_pattern_generator_csr_read),               //                                                .read
		.prbs_pattern_generator_csr_readdata                   (mm_interconnect_0_prbs_pattern_generator_csr_readdata),           //                                                .readdata
		.prbs_pattern_generator_csr_writedata                  (mm_interconnect_0_prbs_pattern_generator_csr_writedata),          //                                                .writedata
		.prbs_pattern_generator_csr_byteenable                 (mm_interconnect_0_prbs_pattern_generator_csr_byteenable),         //                                                .byteenable
		.status_mon_0_slv_address                              (mm_interconnect_0_status_mon_0_slv_address),                      //                                status_mon_0_slv.address
		.status_mon_0_slv_write                                (mm_interconnect_0_status_mon_0_slv_write),                        //                                                .write
		.status_mon_0_slv_read                                 (mm_interconnect_0_status_mon_0_slv_read),                         //                                                .read
		.status_mon_0_slv_readdata                             (mm_interconnect_0_status_mon_0_slv_readdata),                     //                                                .readdata
		.status_mon_0_slv_writedata                            (mm_interconnect_0_status_mon_0_slv_writedata),                    //                                                .writedata
		.status_mon_0_slv_chipselect                           (mm_interconnect_0_status_mon_0_slv_chipselect),                   //                                                .chipselect
		.timer_0_s1_address                                    (mm_interconnect_0_timer_0_s1_address),                            //                                      timer_0_s1.address
		.timer_0_s1_write                                      (mm_interconnect_0_timer_0_s1_write),                              //                                                .write
		.timer_0_s1_readdata                                   (mm_interconnect_0_timer_0_s1_readdata),                           //                                                .readdata
		.timer_0_s1_writedata                                  (mm_interconnect_0_timer_0_s1_writedata),                          //                                                .writedata
		.timer_0_s1_chipselect                                 (mm_interconnect_0_timer_0_s1_chipselect)                          //                                                .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_0_reset_n),                   // reset_in0.reset
		.clk            (clk_0_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_0_reset_n),                   // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_0_clk),                          //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

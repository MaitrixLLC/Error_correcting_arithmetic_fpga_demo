
module global_clk_1 (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
